
module enumerate ( prm, enm );
  input [47:0] prm;
  output [14:0] enm;
  wire   n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364;

  CKND2D0 U84 ( .A1(n321), .A2(prm[0]), .ZN(n70) );
  MAOI222D0 U85 ( .A(n185), .B(prm[19]), .C(n70), .ZN(n71) );
  MAOI222D0 U86 ( .A(n324), .B(prm[2]), .C(n71), .ZN(n72) );
  CKND0 U87 ( .I(n72), .ZN(n73) );
  MAOI222D0 U88 ( .A(prm[3]), .B(n310), .C(n73), .ZN(n74) );
  MAOI222D0 U89 ( .A(prm[22]), .B(n202), .C(n74), .ZN(n75) );
  MAOI222D0 U90 ( .A(n312), .B(prm[5]), .C(n75), .ZN(n204) );
  NR2D0 U91 ( .A1(n292), .A2(prm[18]), .ZN(n76) );
  MAOI222D0 U92 ( .A(prm[7]), .B(n275), .C(n76), .ZN(n77) );
  IAO21D0 U93 ( .A1(prm[20]), .A2(n77), .B(prm[8]), .ZN(n78) );
  MAOI222D0 U94 ( .A(prm[21]), .B(n78), .C(n297), .ZN(n79) );
  OAI211D0 U95 ( .A1(n297), .A2(prm[21]), .B(prm[20]), .C(n77), .ZN(n80) );
  CKND2D0 U96 ( .A1(n79), .A2(n80), .ZN(n81) );
  MAOI222D0 U97 ( .A(n301), .B(prm[22]), .C(n81), .ZN(n82) );
  MAOI222D0 U98 ( .A(n312), .B(prm[11]), .C(n82), .ZN(n278) );
  CKND0 U99 ( .I(prm[28]), .ZN(n83) );
  CKND0 U100 ( .I(prm[26]), .ZN(n84) );
  MAOI222D0 U101 ( .A(prm[25]), .B(n323), .C(n223), .ZN(n85) );
  MAOI222D0 U102 ( .A(prm[32]), .B(n84), .C(n85), .ZN(n86) );
  MAOI222D0 U103 ( .A(n326), .B(prm[27]), .C(n86), .ZN(n87) );
  MAOI222D0 U104 ( .A(prm[34]), .B(n83), .C(n87), .ZN(n88) );
  MAOI222D0 U105 ( .A(n331), .B(prm[29]), .C(n88), .ZN(n89) );
  MAOI222D0 U106 ( .A(prm[38]), .B(n221), .C(n84), .ZN(n90) );
  NR2D0 U107 ( .A1(prm[39]), .A2(n316), .ZN(n91) );
  OAI222D0 U108 ( .A1(n90), .A2(n91), .B1(prm[28]), .B2(n311), .C1(n245), .C2(
        prm[27]), .ZN(n92) );
  OAI21D0 U109 ( .A1(prm[40]), .A2(n83), .B(n92), .ZN(n93) );
  MAOI222D0 U110 ( .A(prm[29]), .B(n303), .C(n93), .ZN(n94) );
  MAOI222D0 U111 ( .A(prm[44]), .B(n219), .C(n84), .ZN(n95) );
  NR2D0 U112 ( .A1(prm[45]), .A2(n316), .ZN(n96) );
  OAI222D0 U113 ( .A1(n95), .A2(n96), .B1(prm[28]), .B2(n308), .C1(n286), .C2(
        prm[27]), .ZN(n97) );
  OAI21D0 U114 ( .A1(prm[46]), .A2(n83), .B(n97), .ZN(n98) );
  MAOI222D0 U115 ( .A(prm[29]), .B(n291), .C(n98), .ZN(n99) );
  MAOI222D0 U116 ( .A(n89), .B(n94), .C(n99), .ZN(n100) );
  CKND0 U117 ( .I(n100), .ZN(n224) );
  XOR3D0 U118 ( .A1(n89), .A2(n94), .A3(n99), .Z(n225) );
  NR2D0 U119 ( .A1(n193), .A2(prm[24]), .ZN(n101) );
  MAOI222D0 U120 ( .A(prm[1]), .B(n314), .C(n101), .ZN(n102) );
  IAO21D0 U121 ( .A1(prm[26]), .A2(n102), .B(prm[2]), .ZN(n103) );
  MAOI222D0 U122 ( .A(prm[27]), .B(n103), .C(n197), .ZN(n104) );
  OAI211D0 U123 ( .A1(n197), .A2(prm[27]), .B(prm[26]), .C(n102), .ZN(n105) );
  CKND2D0 U124 ( .A1(n104), .A2(n105), .ZN(n106) );
  MAOI222D0 U125 ( .A(n202), .B(prm[28]), .C(n106), .ZN(n107) );
  MAOI222D0 U126 ( .A(n320), .B(prm[5]), .C(n107), .ZN(n205) );
  NR2D0 U127 ( .A1(n292), .A2(prm[12]), .ZN(n108) );
  MAOI222D0 U128 ( .A(prm[7]), .B(n273), .C(n108), .ZN(n109) );
  OAI211D0 U129 ( .A1(n297), .A2(prm[15]), .B(prm[14]), .C(n109), .ZN(n110) );
  IAO21D0 U130 ( .A1(prm[14]), .A2(n109), .B(prm[8]), .ZN(n111) );
  MAOI222D0 U131 ( .A(n297), .B(n111), .C(prm[15]), .ZN(n112) );
  CKND2D0 U132 ( .A1(n112), .A2(n110), .ZN(n113) );
  MAOI222D0 U133 ( .A(prm[16]), .B(n301), .C(n113), .ZN(n114) );
  MAOI222D0 U134 ( .A(n274), .B(prm[11]), .C(n114), .ZN(n279) );
  NR2D0 U135 ( .A1(prm[36]), .A2(n321), .ZN(n115) );
  MAOI222D0 U136 ( .A(n309), .B(prm[19]), .C(n115), .ZN(n116) );
  MAOI222D0 U137 ( .A(n324), .B(prm[38]), .C(n116), .ZN(n117) );
  CKND0 U138 ( .I(n117), .ZN(n118) );
  MAOI222D0 U139 ( .A(prm[39]), .B(n310), .C(n118), .ZN(n119) );
  MAOI222D0 U140 ( .A(prm[22]), .B(n311), .C(n119), .ZN(n120) );
  MAOI222D0 U141 ( .A(prm[41]), .B(n312), .C(n120), .ZN(n351) );
  NR2D0 U142 ( .A1(prm[42]), .A2(n226), .ZN(n121) );
  MAOI222D0 U143 ( .A(prm[31]), .B(n307), .C(n121), .ZN(n122) );
  MAOI222D0 U144 ( .A(n227), .B(prm[44]), .C(n122), .ZN(n123) );
  CKND0 U145 ( .I(n123), .ZN(n124) );
  MAOI222D0 U146 ( .A(prm[45]), .B(n326), .C(n124), .ZN(n125) );
  MAOI222D0 U147 ( .A(prm[34]), .B(n308), .C(n125), .ZN(n126) );
  MAOI222D0 U148 ( .A(prm[47]), .B(n331), .C(n126), .ZN(n266) );
  NR2D0 U149 ( .A1(n292), .A2(prm[24]), .ZN(n127) );
  MAOI222D0 U150 ( .A(prm[7]), .B(n314), .C(n127), .ZN(n128) );
  IAO21D0 U151 ( .A1(prm[26]), .A2(n128), .B(prm[8]), .ZN(n129) );
  OAI211D0 U152 ( .A1(n297), .A2(prm[27]), .B(prm[26]), .C(n128), .ZN(n130) );
  MAOI222D0 U153 ( .A(prm[27]), .B(n129), .C(n297), .ZN(n131) );
  CKND2D0 U154 ( .A1(n131), .A2(n130), .ZN(n132) );
  MAOI222D0 U155 ( .A(n301), .B(prm[28]), .C(n132), .ZN(n133) );
  MAOI222D0 U156 ( .A(n320), .B(prm[11]), .C(n133), .ZN(n277) );
  NR2D0 U157 ( .A1(prm[42]), .A2(n321), .ZN(n134) );
  MAOI222D0 U158 ( .A(n307), .B(prm[19]), .C(n134), .ZN(n135) );
  MAOI222D0 U159 ( .A(n324), .B(prm[44]), .C(n135), .ZN(n136) );
  CKND0 U160 ( .I(n136), .ZN(n137) );
  MAOI222D0 U161 ( .A(prm[45]), .B(n310), .C(n137), .ZN(n138) );
  MAOI222D0 U162 ( .A(prm[22]), .B(n308), .C(n138), .ZN(n139) );
  MAOI222D0 U163 ( .A(prm[47]), .B(n312), .C(n139), .ZN(n352) );
  NR2D0 U164 ( .A1(prm[36]), .A2(n226), .ZN(n140) );
  MAOI222D0 U165 ( .A(prm[31]), .B(n309), .C(n140), .ZN(n141) );
  MAOI222D0 U166 ( .A(n227), .B(prm[38]), .C(n141), .ZN(n142) );
  CKND0 U167 ( .I(n142), .ZN(n143) );
  MAOI222D0 U168 ( .A(prm[39]), .B(n326), .C(n143), .ZN(n144) );
  MAOI222D0 U169 ( .A(prm[34]), .B(n311), .C(n144), .ZN(n145) );
  MAOI222D0 U170 ( .A(prm[41]), .B(n331), .C(n145), .ZN(n265) );
  NR2D0 U171 ( .A1(n292), .A2(prm[30]), .ZN(n146) );
  MAOI222D0 U172 ( .A(prm[7]), .B(n323), .C(n146), .ZN(n147) );
  IAO21D0 U173 ( .A1(prm[32]), .A2(n147), .B(prm[8]), .ZN(n148) );
  OAI211D0 U174 ( .A1(n297), .A2(prm[33]), .B(prm[32]), .C(n147), .ZN(n149) );
  MAOI222D0 U175 ( .A(prm[33]), .B(n148), .C(n297), .ZN(n150) );
  CKND2D0 U176 ( .A1(n150), .A2(n149), .ZN(n151) );
  MAOI222D0 U177 ( .A(n301), .B(prm[34]), .C(n151), .ZN(n152) );
  MAOI222D0 U178 ( .A(n331), .B(prm[11]), .C(n152), .ZN(n276) );
  AOI22D0 U179 ( .A1(n211), .A2(n212), .B1(n213), .B2(n217), .ZN(n153) );
  OAI21D0 U180 ( .A1(n213), .A2(n217), .B(n153), .ZN(n268) );
  CKND0 U181 ( .I(prm[42]), .ZN(n154) );
  OAI211D0 U182 ( .A1(prm[37]), .A2(n307), .B(prm[36]), .C(n154), .ZN(n155) );
  OAI21D0 U183 ( .A1(prm[43]), .A2(n309), .B(n155), .ZN(n156) );
  AOI211D0 U184 ( .A1(prm[39]), .A2(n286), .B(prm[38]), .C(n156), .ZN(n157) );
  IOA21D0 U185 ( .A1(prm[38]), .A2(n156), .B(prm[44]), .ZN(n158) );
  MAOI222D0 U186 ( .A(n286), .B(prm[39]), .C(n158), .ZN(n159) );
  NR2D0 U187 ( .A1(n157), .A2(n159), .ZN(n160) );
  MAOI222D0 U188 ( .A(prm[40]), .B(n308), .C(n160), .ZN(n161) );
  MAOI222D0 U189 ( .A(prm[47]), .B(n303), .C(n161), .ZN(enm[14]) );
  CKND0 U190 ( .I(n269), .ZN(n214) );
  CKND0 U191 ( .I(n213), .ZN(n216) );
  CKND2D0 U192 ( .A1(n346), .A2(n267), .ZN(enm[13]) );
  CKND2D0 U193 ( .A1(n345), .A2(n344), .ZN(n267) );
  CKND0 U194 ( .I(n225), .ZN(enm[11]) );
  CKND0 U195 ( .I(n224), .ZN(enm[10]) );
  CKND0 U196 ( .I(prm[24]), .ZN(n222) );
  CKND2D0 U197 ( .A1(n360), .A2(n359), .ZN(n358) );
  CKND0 U198 ( .I(n350), .ZN(enm[7]) );
  CKND0 U199 ( .I(n343), .ZN(n344) );
  CKND0 U200 ( .I(n342), .ZN(n345) );
  CKND0 U201 ( .I(prm[12]), .ZN(n254) );
  CKND0 U202 ( .I(prm[14]), .ZN(n257) );
  CKND0 U203 ( .I(n357), .ZN(n363) );
  CKND0 U204 ( .I(n336), .ZN(n337) );
  CKND0 U205 ( .I(prm[27]), .ZN(n316) );
  CKND0 U206 ( .I(prm[22]), .ZN(n329) );
  CKND0 U207 ( .I(n362), .ZN(n338) );
  CKND2D0 U208 ( .A1(n352), .A2(n351), .ZN(n362) );
  CKND0 U209 ( .I(prm[40]), .ZN(n311) );
  CKND0 U210 ( .I(prm[37]), .ZN(n309) );
  CKND0 U211 ( .I(prm[46]), .ZN(n308) );
  CKND0 U212 ( .I(prm[8]), .ZN(n294) );
  CKND0 U213 ( .I(n332), .ZN(n281) );
  CKND0 U214 ( .I(prm[19]), .ZN(n275) );
  CKND0 U215 ( .I(prm[31]), .ZN(n323) );
  CKND0 U216 ( .I(prm[6]), .ZN(n292) );
  OR2D0 U217 ( .A1(n204), .A2(n205), .Z(n217) );
  CKND2D0 U218 ( .A1(n173), .A2(n172), .ZN(n174) );
  CKND2D0 U219 ( .A1(prm[3]), .A2(n326), .ZN(n172) );
  CKND0 U220 ( .I(prm[32]), .ZN(n227) );
  CKND2D0 U221 ( .A1(prm[0]), .A2(n226), .ZN(n170) );
  CKND0 U222 ( .I(prm[30]), .ZN(n226) );
  CKND0 U223 ( .I(prm[33]), .ZN(n326) );
  CKND2D0 U224 ( .A1(n185), .A2(n193), .ZN(n165) );
  CKND0 U225 ( .I(prm[39]), .ZN(n245) );
  CKND2D0 U226 ( .A1(prm[1]), .A2(prm[0]), .ZN(n162) );
  CKND0 U227 ( .I(prm[20]), .ZN(n324) );
  CKND0 U228 ( .I(prm[18]), .ZN(n321) );
  CKND0 U229 ( .I(prm[21]), .ZN(n310) );
  CKND0 U230 ( .I(prm[25]), .ZN(n314) );
  CKND0 U231 ( .I(prm[29]), .ZN(n320) );
  CKND0 U232 ( .I(prm[13]), .ZN(n273) );
  CKND0 U233 ( .I(prm[15]), .ZN(n248) );
  CKND0 U234 ( .I(prm[16]), .ZN(n260) );
  CKND0 U235 ( .I(prm[17]), .ZN(n274) );
  CKND0 U236 ( .I(prm[45]), .ZN(n286) );
  CKND0 U237 ( .I(prm[1]), .ZN(n185) );
  CKND0 U238 ( .I(prm[43]), .ZN(n307) );
  CKND0 U239 ( .I(prm[47]), .ZN(n291) );
  CKND0 U240 ( .I(prm[3]), .ZN(n197) );
  CKND0 U241 ( .I(prm[2]), .ZN(n195) );
  CKND0 U242 ( .I(prm[0]), .ZN(n193) );
  CKND0 U243 ( .I(prm[7]), .ZN(n282) );
  CKND0 U244 ( .I(prm[9]), .ZN(n297) );
  CKND0 U245 ( .I(prm[10]), .ZN(n301) );
  CKND0 U246 ( .I(prm[4]), .ZN(n202) );
  CKND0 U247 ( .I(prm[11]), .ZN(n184) );
  INVD1 U248 ( .I(prm[35]), .ZN(n331) );
  OAI21D1 U249 ( .A1(n217), .A2(n216), .B(n215), .ZN(enm[0]) );
  MAOI222D1 U250 ( .A(n270), .B(n214), .C(n268), .ZN(n215) );
  IOA21D1 U251 ( .A1(n266), .A2(n265), .B(n267), .ZN(enm[12]) );
  NR2D1 U252 ( .A1(n222), .A2(prm[30]), .ZN(n223) );
  MAOI222D1 U253 ( .A(prm[25]), .B(n309), .C(n220), .ZN(n221) );
  NR2D1 U254 ( .A1(n222), .A2(prm[36]), .ZN(n220) );
  MAOI222D1 U255 ( .A(prm[25]), .B(n307), .C(n218), .ZN(n219) );
  NR2D1 U256 ( .A1(n222), .A2(prm[42]), .ZN(n218) );
  OAI31D1 U257 ( .A1(n364), .A2(n363), .A3(n362), .B(n361), .ZN(enm[9]) );
  OAI21D1 U258 ( .A1(n360), .A2(n359), .B(n358), .ZN(n361) );
  OAI211D1 U259 ( .A1(n357), .A2(n362), .B(n358), .C(n356), .ZN(enm[8]) );
  OAI21D1 U260 ( .A1(n362), .A2(n355), .B(n357), .ZN(n356) );
  CKXOR2D1 U261 ( .A1(n354), .A2(n353), .Z(n359) );
  CKXOR2D1 U262 ( .A1(n352), .A2(n351), .Z(n360) );
  AOI32D1 U263 ( .A1(n346), .A2(n345), .A3(n344), .B1(n343), .B2(n342), .ZN(
        enm[6]) );
  MAOI222D1 U264 ( .A(prm[17]), .B(n331), .C(n261), .ZN(n347) );
  MAOI222D1 U265 ( .A(prm[34]), .B(n260), .C(n259), .ZN(n261) );
  MAOI222D1 U266 ( .A(prm[15]), .B(n258), .C(n326), .ZN(n259) );
  MAOI222D1 U267 ( .A(prm[32]), .B(n257), .C(n256), .ZN(n258) );
  MAOI222D1 U268 ( .A(prm[13]), .B(n323), .C(n255), .ZN(n256) );
  NR2D1 U269 ( .A1(n254), .A2(prm[30]), .ZN(n255) );
  MAOI222D1 U270 ( .A(prm[17]), .B(n303), .C(n253), .ZN(n348) );
  OAI22D1 U271 ( .A1(prm[40]), .A2(n260), .B1(n252), .B2(n251), .ZN(n253) );
  NR2D1 U272 ( .A1(n250), .A2(n249), .ZN(n251) );
  NR2D1 U273 ( .A1(prm[39]), .A2(n248), .ZN(n249) );
  MAOI222D1 U274 ( .A(n247), .B(prm[38]), .C(n257), .ZN(n250) );
  MAOI222D1 U275 ( .A(prm[13]), .B(n309), .C(n246), .ZN(n247) );
  NR2D1 U276 ( .A1(n254), .A2(prm[36]), .ZN(n246) );
  OAI22D1 U277 ( .A1(prm[16]), .A2(n311), .B1(prm[15]), .B2(n245), .ZN(n252)
         );
  MAOI222D1 U278 ( .A(prm[17]), .B(n320), .C(n244), .ZN(n262) );
  MAOI222D1 U279 ( .A(prm[28]), .B(n260), .C(n243), .ZN(n244) );
  MAOI222D1 U280 ( .A(prm[15]), .B(n242), .C(n316), .ZN(n243) );
  MAOI222D1 U281 ( .A(prm[26]), .B(n257), .C(n241), .ZN(n242) );
  MAOI222D1 U282 ( .A(prm[13]), .B(n314), .C(n240), .ZN(n241) );
  NR2D1 U283 ( .A1(n254), .A2(prm[24]), .ZN(n240) );
  MAOI222D1 U284 ( .A(prm[17]), .B(n291), .C(n239), .ZN(n263) );
  OAI22D1 U285 ( .A1(prm[46]), .A2(n260), .B1(n238), .B2(n237), .ZN(n239) );
  NR2D1 U286 ( .A1(n236), .A2(n235), .ZN(n237) );
  NR2D1 U287 ( .A1(prm[45]), .A2(n248), .ZN(n235) );
  MAOI222D1 U288 ( .A(n234), .B(prm[44]), .C(n257), .ZN(n236) );
  MAOI222D1 U289 ( .A(prm[13]), .B(n307), .C(n233), .ZN(n234) );
  NR2D1 U290 ( .A1(n254), .A2(prm[42]), .ZN(n233) );
  OAI22D1 U291 ( .A1(prm[16]), .A2(n308), .B1(prm[15]), .B2(n286), .ZN(n238)
         );
  MAOI222D1 U292 ( .A(prm[17]), .B(n312), .C(n232), .ZN(n264) );
  MAOI222D1 U293 ( .A(prm[22]), .B(n260), .C(n231), .ZN(n232) );
  MAOI222D1 U294 ( .A(prm[15]), .B(n230), .C(n310), .ZN(n231) );
  MAOI222D1 U295 ( .A(prm[20]), .B(n257), .C(n229), .ZN(n230) );
  MAOI222D1 U296 ( .A(prm[13]), .B(n275), .C(n228), .ZN(n229) );
  NR2D1 U297 ( .A1(n254), .A2(prm[18]), .ZN(n228) );
  XNR2D1 U298 ( .A1(n266), .A2(n265), .ZN(n346) );
  OAI21D1 U299 ( .A1(n362), .A2(n363), .B(n364), .ZN(enm[5]) );
  AO21D1 U300 ( .A1(n357), .A2(n338), .B(n355), .Z(enm[4]) );
  OAI21D1 U301 ( .A1(n335), .A2(n336), .B(n334), .ZN(enm[3]) );
  AOI22D1 U302 ( .A1(n338), .A2(n357), .B1(n333), .B2(n332), .ZN(n334) );
  NR2D1 U303 ( .A1(n353), .A2(n354), .ZN(n357) );
  MAOI222D1 U304 ( .A(prm[23]), .B(n331), .C(n330), .ZN(n354) );
  MAOI222D1 U305 ( .A(prm[34]), .B(n329), .C(n328), .ZN(n330) );
  MAOI222D1 U306 ( .A(n327), .B(prm[21]), .C(n326), .ZN(n328) );
  MAOI222D1 U307 ( .A(prm[32]), .B(n325), .C(n324), .ZN(n327) );
  MAOI222D1 U308 ( .A(prm[19]), .B(n323), .C(n322), .ZN(n325) );
  NR2D1 U309 ( .A1(n321), .A2(prm[30]), .ZN(n322) );
  MAOI222D1 U310 ( .A(prm[23]), .B(n320), .C(n319), .ZN(n353) );
  MAOI222D1 U311 ( .A(prm[28]), .B(n329), .C(n318), .ZN(n319) );
  MAOI222D1 U312 ( .A(n317), .B(prm[21]), .C(n316), .ZN(n318) );
  MAOI222D1 U313 ( .A(prm[26]), .B(n315), .C(n324), .ZN(n317) );
  MAOI222D1 U314 ( .A(prm[19]), .B(n314), .C(n313), .ZN(n315) );
  NR2D1 U315 ( .A1(n321), .A2(prm[24]), .ZN(n313) );
  AO21D1 U316 ( .A1(n306), .A2(n305), .B(n304), .Z(n339) );
  MAOI222D1 U317 ( .A(prm[11]), .B(n303), .C(n302), .ZN(n340) );
  MAOI222D1 U318 ( .A(prm[40]), .B(n301), .C(n300), .ZN(n302) );
  OAI21D1 U319 ( .A1(prm[8]), .A2(n299), .B(n298), .ZN(n300) );
  AOI22D1 U320 ( .A1(prm[39]), .A2(n297), .B1(n296), .B2(n295), .ZN(n298) );
  MAOI222D1 U321 ( .A(prm[7]), .B(n309), .C(n293), .ZN(n296) );
  NR2D1 U322 ( .A1(n292), .A2(prm[36]), .ZN(n293) );
  OAI21D1 U323 ( .A1(prm[39]), .A2(n297), .B(prm[38]), .ZN(n299) );
  MAOI222D1 U324 ( .A(prm[11]), .B(n291), .C(n290), .ZN(n341) );
  OAI22D1 U325 ( .A1(prm[46]), .A2(n301), .B1(n289), .B2(n288), .ZN(n290) );
  OAI22D1 U326 ( .A1(prm[10]), .A2(n308), .B1(prm[8]), .B2(n287), .ZN(n288) );
  OAI21D1 U327 ( .A1(prm[45]), .A2(n297), .B(prm[44]), .ZN(n287) );
  OAI22D1 U328 ( .A1(prm[9]), .A2(n286), .B1(n285), .B2(n284), .ZN(n289) );
  OAI22D1 U329 ( .A1(prm[45]), .A2(n297), .B1(prm[44]), .B2(n294), .ZN(n284)
         );
  OAI32D1 U330 ( .A1(n283), .A2(n292), .A3(prm[42]), .B1(prm[43]), .B2(n282), 
        .ZN(n285) );
  NR2D1 U331 ( .A1(prm[7]), .A2(n307), .ZN(n283) );
  AOI211D1 U332 ( .A1(n333), .A2(n281), .B(n304), .C(n280), .ZN(n335) );
  NR2D1 U333 ( .A1(n333), .A2(n281), .ZN(n280) );
  NR2D1 U334 ( .A1(n306), .A2(n305), .ZN(n304) );
  XNR2D1 U335 ( .A1(n279), .A2(n278), .ZN(n305) );
  XNR2D1 U336 ( .A1(n277), .A2(n276), .ZN(n306) );
  NR2D1 U337 ( .A1(n279), .A2(n278), .ZN(n332) );
  NR2D1 U338 ( .A1(n277), .A2(n276), .ZN(n333) );
  AOI21D1 U339 ( .A1(n272), .A2(n271), .B(n270), .ZN(enm[2]) );
  XNR3D1 U340 ( .A1(n270), .A2(n269), .A3(n268), .ZN(enm[1]) );
  NR2D1 U341 ( .A1(n207), .A2(n206), .ZN(n213) );
  NR2D1 U342 ( .A1(n272), .A2(n271), .ZN(n270) );
  XNR2D1 U343 ( .A1(n212), .A2(n211), .ZN(n271) );
  CKXOR2D1 U344 ( .A1(n207), .A2(n206), .Z(n211) );
  MAOI222D1 U345 ( .A(prm[5]), .B(n331), .C(n176), .ZN(n206) );
  MAOI222D1 U346 ( .A(prm[34]), .B(n202), .C(n175), .ZN(n176) );
  OAI21D1 U347 ( .A1(prm[3]), .A2(n326), .B(n174), .ZN(n175) );
  MAOI222D1 U348 ( .A(prm[2]), .B(n171), .C(n227), .ZN(n173) );
  MAOI222D1 U349 ( .A(prm[31]), .B(n170), .C(n185), .ZN(n171) );
  MAOI222D1 U350 ( .A(prm[5]), .B(n303), .C(n169), .ZN(n207) );
  MAOI222D1 U351 ( .A(prm[40]), .B(n202), .C(n168), .ZN(n169) );
  AOI32D1 U352 ( .A1(n167), .A2(n166), .A3(n165), .B1(n164), .B2(n166), .ZN(
        n168) );
  OAI22D1 U353 ( .A1(prm[39]), .A2(n197), .B1(prm[38]), .B2(n195), .ZN(n164)
         );
  AOI22D1 U354 ( .A1(prm[39]), .A2(n197), .B1(prm[38]), .B2(n163), .ZN(n166)
         );
  AOI21D1 U355 ( .A1(prm[3]), .A2(n245), .B(prm[2]), .ZN(n163) );
  INVD1 U356 ( .I(prm[41]), .ZN(n303) );
  CKXOR2D1 U357 ( .A1(n205), .A2(n204), .Z(n212) );
  INVD1 U358 ( .I(prm[23]), .ZN(n312) );
  MAOI222D1 U359 ( .A(prm[5]), .B(n274), .C(n203), .ZN(n208) );
  OAI22D1 U360 ( .A1(prm[16]), .A2(n202), .B1(n201), .B2(n200), .ZN(n203) );
  NR2D1 U361 ( .A1(n199), .A2(n198), .ZN(n200) );
  NR2D1 U362 ( .A1(prm[15]), .A2(n197), .ZN(n198) );
  MAOI222D1 U363 ( .A(n196), .B(prm[14]), .C(n195), .ZN(n199) );
  MAOI222D1 U364 ( .A(prm[1]), .B(n273), .C(n194), .ZN(n196) );
  NR2D1 U365 ( .A1(n193), .A2(prm[12]), .ZN(n194) );
  OAI22D1 U366 ( .A1(prm[4]), .A2(n260), .B1(prm[3]), .B2(n248), .ZN(n201) );
  MAOI222D1 U367 ( .A(prm[5]), .B(n291), .C(n192), .ZN(n209) );
  MAOI222D1 U368 ( .A(prm[46]), .B(n202), .C(n191), .ZN(n192) );
  OAI21D1 U369 ( .A1(n190), .A2(n189), .B(n188), .ZN(n191) );
  AOI22D1 U370 ( .A1(prm[45]), .A2(n197), .B1(prm[44]), .B2(n187), .ZN(n188)
         );
  AOI21D1 U371 ( .A1(prm[3]), .A2(n286), .B(prm[2]), .ZN(n187) );
  OAI22D1 U372 ( .A1(prm[45]), .A2(n197), .B1(prm[44]), .B2(n195), .ZN(n189)
         );
  OAI32D1 U373 ( .A1(n186), .A2(n193), .A3(prm[42]), .B1(prm[43]), .B2(n185), 
        .ZN(n190) );
  NR2D1 U374 ( .A1(prm[1]), .A2(n307), .ZN(n186) );
  MAOI222D1 U375 ( .A(prm[5]), .B(n184), .C(n183), .ZN(n210) );
  OAI22D1 U376 ( .A1(prm[10]), .A2(n202), .B1(n182), .B2(n181), .ZN(n183) );
  NR2D1 U377 ( .A1(n180), .A2(n179), .ZN(n181) );
  NR2D1 U378 ( .A1(prm[9]), .A2(n197), .ZN(n179) );
  MAOI222D1 U379 ( .A(n178), .B(prm[8]), .C(n195), .ZN(n180) );
  MAOI222D1 U380 ( .A(prm[1]), .B(n282), .C(n177), .ZN(n178) );
  NR2D1 U381 ( .A1(n193), .A2(prm[6]), .ZN(n177) );
  OAI22D1 U382 ( .A1(prm[4]), .A2(n301), .B1(prm[3]), .B2(n297), .ZN(n182) );
  OAI222D0 U383 ( .A1(prm[37]), .A2(n185), .B1(prm[37]), .B2(prm[36]), .C1(
        prm[36]), .C2(n162), .ZN(n167) );
  FA1D0 U384 ( .A(n210), .B(n209), .CI(n208), .CO(n269), .S(n272) );
  FA1D0 U385 ( .A(n264), .B(n263), .CI(n262), .CO(n343), .S(n349) );
  OA22D0 U386 ( .A1(n297), .A2(prm[39]), .B1(n294), .B2(prm[38]), .Z(n295) );
  MUX2ND0 U387 ( .I0(n337), .I1(n336), .S(n335), .ZN(n355) );
  FA1D0 U388 ( .A(n341), .B(n340), .CI(n339), .CO(n336), .S(n364) );
  FA1D0 U389 ( .A(n349), .B(n348), .CI(n347), .CO(n342), .S(n350) );
endmodule

