
module enumerate ( prm, enm );
  input [41:0] prm;
  output [11:0] enm;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261;

  CKND0 U62 ( .I(prm[11]), .ZN(n51) );
  CKND2D0 U63 ( .A1(n175), .A2(prm[0]), .ZN(n52) );
  MAOI222D0 U64 ( .A(n111), .B(prm[7]), .C(n52), .ZN(n53) );
  MAOI222D0 U65 ( .A(n178), .B(prm[2]), .C(n53), .ZN(n54) );
  CKND0 U66 ( .I(n54), .ZN(n55) );
  MAOI222D0 U67 ( .A(prm[3]), .B(n153), .C(n55), .ZN(n56) );
  MAOI222D0 U68 ( .A(prm[10]), .B(n118), .C(n56), .ZN(n57) );
  MAOI222D0 U69 ( .A(prm[5]), .B(n51), .C(n57), .ZN(n100) );
  CKND2D0 U70 ( .A1(n133), .A2(prm[0]), .ZN(n58) );
  MAOI222D0 U71 ( .A(prm[13]), .B(n111), .C(n58), .ZN(n59) );
  MAOI222D0 U72 ( .A(n136), .B(prm[2]), .C(n59), .ZN(n60) );
  MAOI222D0 U73 ( .A(prm[3]), .B(n61), .C(n62), .ZN(n63) );
  MAOI222D0 U74 ( .A(prm[16]), .B(n118), .C(n63), .ZN(n64) );
  MAOI222D0 U75 ( .A(n166), .B(prm[5]), .C(n64), .ZN(n99) );
  CKND0 U76 ( .I(n60), .ZN(n61) );
  CKND0 U77 ( .I(prm[15]), .ZN(n62) );
  CKND2D0 U78 ( .A1(prm[0]), .A2(n191), .ZN(n65) );
  MAOI222D0 U79 ( .A(prm[25]), .B(n111), .C(n65), .ZN(n66) );
  MAOI222D0 U80 ( .A(n192), .B(prm[2]), .C(n66), .ZN(n67) );
  CKND0 U81 ( .I(n67), .ZN(n68) );
  MAOI222D0 U82 ( .A(prm[3]), .B(n248), .C(n68), .ZN(n69) );
  MAOI222D0 U83 ( .A(n118), .B(prm[28]), .C(n69), .ZN(n70) );
  MAOI222D0 U84 ( .A(n253), .B(prm[5]), .C(n70), .ZN(n97) );
  NR2D0 U85 ( .A1(prm[36]), .A2(n133), .ZN(n71) );
  MAOI222D0 U86 ( .A(n226), .B(prm[13]), .C(n71), .ZN(n72) );
  MAOI222D0 U87 ( .A(n136), .B(prm[38]), .C(n72), .ZN(n73) );
  CKND0 U88 ( .I(n73), .ZN(n74) );
  MAOI222D0 U89 ( .A(prm[39]), .B(n162), .C(n74), .ZN(n75) );
  MAOI222D0 U90 ( .A(prm[16]), .B(n224), .C(n75), .ZN(n76) );
  MAOI222D0 U91 ( .A(prm[41]), .B(n166), .C(n76), .ZN(n209) );
  CKND2D0 U92 ( .A1(prm[0]), .A2(n243), .ZN(n77) );
  MAOI222D0 U93 ( .A(n111), .B(prm[19]), .C(n77), .ZN(n78) );
  MAOI222D0 U94 ( .A(n247), .B(prm[2]), .C(n78), .ZN(n79) );
  CKND0 U95 ( .I(n79), .ZN(n80) );
  MAOI222D0 U96 ( .A(prm[3]), .B(n228), .C(n80), .ZN(n81) );
  MAOI222D0 U97 ( .A(prm[22]), .B(n118), .C(n81), .ZN(n82) );
  MAOI222D0 U98 ( .A(n150), .B(prm[5]), .C(n82), .ZN(n98) );
  NR2D0 U99 ( .A1(prm[36]), .A2(n191), .ZN(n83) );
  MAOI222D0 U100 ( .A(prm[25]), .B(n226), .C(n83), .ZN(n84) );
  MAOI222D0 U101 ( .A(n192), .B(prm[38]), .C(n84), .ZN(n85) );
  CKND0 U102 ( .I(n85), .ZN(n86) );
  MAOI222D0 U103 ( .A(n248), .B(prm[39]), .C(n86), .ZN(n87) );
  MAOI222D0 U104 ( .A(prm[28]), .B(n224), .C(n87), .ZN(n88) );
  MAOI222D0 U105 ( .A(prm[41]), .B(n253), .C(n88), .ZN(n260) );
  CKND2D0 U106 ( .A1(n259), .A2(n204), .ZN(enm[10]) );
  CKND2D0 U107 ( .A1(n202), .A2(n203), .ZN(n259) );
  CKND0 U108 ( .I(n258), .ZN(enm[8]) );
  CKND0 U109 ( .I(n254), .ZN(enm[7]) );
  CKND0 U110 ( .I(prm[22]), .ZN(n251) );
  CKND2D0 U111 ( .A1(prm[38]), .A2(n90), .ZN(n91) );
  CKND2D0 U112 ( .A1(prm[32]), .A2(n92), .ZN(n90) );
  CKND2D0 U113 ( .A1(n218), .A2(n217), .ZN(n216) );
  CKND0 U114 ( .I(n208), .ZN(enm[4]) );
  CKND0 U115 ( .I(n201), .ZN(n202) );
  CKND0 U116 ( .I(n200), .ZN(n203) );
  CKND0 U117 ( .I(prm[31]), .ZN(n236) );
  CKND0 U118 ( .I(prm[10]), .ZN(n181) );
  CKND2D0 U119 ( .A1(prm[24]), .A2(n183), .ZN(n184) );
  CKND0 U120 ( .I(n215), .ZN(n221) );
  CKND0 U121 ( .I(n141), .ZN(n102) );
  CKND0 U122 ( .I(n194), .ZN(n195) );
  CKND0 U123 ( .I(prm[8]), .ZN(n178) );
  CKND0 U124 ( .I(prm[6]), .ZN(n175) );
  CKND0 U125 ( .I(prm[9]), .ZN(n153) );
  CKND0 U126 ( .I(prm[26]), .ZN(n192) );
  CKND0 U127 ( .I(prm[24]), .ZN(n191) );
  CKND0 U128 ( .I(prm[20]), .ZN(n247) );
  CKND0 U129 ( .I(prm[18]), .ZN(n243) );
  CKND2D0 U130 ( .A1(n115), .A2(n114), .ZN(n116) );
  CKND2D0 U131 ( .A1(prm[3]), .A2(n238), .ZN(n114) );
  CKND0 U132 ( .I(prm[1]), .ZN(n111) );
  CKND2D0 U133 ( .A1(prm[0]), .A2(n183), .ZN(n112) );
  CKND0 U134 ( .I(prm[33]), .ZN(n238) );
  CKND0 U135 ( .I(prm[38]), .ZN(n104) );
  CKND0 U136 ( .I(prm[39]), .ZN(n223) );
  CKND0 U137 ( .I(prm[4]), .ZN(n118) );
  CKND0 U138 ( .I(prm[41]), .ZN(n234) );
  CKND0 U139 ( .I(n220), .ZN(n196) );
  CKND2D0 U140 ( .A1(n209), .A2(n210), .ZN(n220) );
  CKND0 U141 ( .I(prm[34]), .ZN(n188) );
  CKND0 U142 ( .I(prm[32]), .ZN(n185) );
  CKND0 U143 ( .I(prm[13]), .ZN(n159) );
  CKND2D0 U144 ( .A1(prm[12]), .A2(n183), .ZN(n123) );
  CKND0 U145 ( .I(prm[30]), .ZN(n183) );
  CKND0 U146 ( .I(prm[17]), .ZN(n166) );
  CKND0 U147 ( .I(prm[40]), .ZN(n224) );
  CKND0 U148 ( .I(prm[37]), .ZN(n226) );
  CKND0 U149 ( .I(prm[15]), .ZN(n162) );
  CKND0 U150 ( .I(prm[27]), .ZN(n248) );
  CKND0 U151 ( .I(prm[25]), .ZN(n245) );
  CKND0 U152 ( .I(prm[21]), .ZN(n228) );
  CKND0 U153 ( .I(prm[14]), .ZN(n136) );
  CKND0 U154 ( .I(prm[12]), .ZN(n133) );
  CKND0 U155 ( .I(prm[19]), .ZN(n145) );
  CKND0 U156 ( .I(prm[16]), .ZN(n139) );
  CKND0 U157 ( .I(prm[23]), .ZN(n150) );
  OAI21D1 U158 ( .A1(n193), .A2(n194), .B(n143), .ZN(enm[0]) );
  AOI22D1 U159 ( .A1(n196), .A2(n215), .B1(n142), .B2(n141), .ZN(n143) );
  IOA21D1 U160 ( .A1(n261), .A2(n260), .B(n259), .ZN(enm[9]) );
  MAOI222D1 U161 ( .A(prm[23]), .B(n253), .C(n252), .ZN(n255) );
  MAOI222D1 U162 ( .A(prm[28]), .B(n251), .C(n250), .ZN(n252) );
  MAOI222D1 U163 ( .A(prm[21]), .B(n249), .C(n248), .ZN(n250) );
  MAOI222D1 U164 ( .A(prm[26]), .B(n247), .C(n246), .ZN(n249) );
  MAOI222D1 U165 ( .A(prm[19]), .B(n245), .C(n244), .ZN(n246) );
  NR2D1 U166 ( .A1(n243), .A2(prm[24]), .ZN(n244) );
  MAOI222D1 U167 ( .A(prm[23]), .B(n242), .C(n241), .ZN(n256) );
  MAOI222D1 U168 ( .A(prm[34]), .B(n251), .C(n240), .ZN(n241) );
  MAOI222D1 U169 ( .A(prm[21]), .B(n239), .C(n238), .ZN(n240) );
  MAOI222D1 U170 ( .A(prm[32]), .B(n247), .C(n237), .ZN(n239) );
  MAOI222D1 U171 ( .A(prm[19]), .B(n236), .C(n235), .ZN(n237) );
  NR2D1 U172 ( .A1(n243), .A2(prm[30]), .ZN(n235) );
  MAOI222D1 U173 ( .A(prm[23]), .B(n234), .C(n233), .ZN(n257) );
  OAI22D1 U174 ( .A1(prm[40]), .A2(n251), .B1(n232), .B2(n231), .ZN(n233) );
  NR2D1 U175 ( .A1(n230), .A2(n229), .ZN(n231) );
  NR2D1 U176 ( .A1(prm[39]), .A2(n228), .ZN(n229) );
  MAOI222D1 U177 ( .A(n227), .B(prm[38]), .C(n247), .ZN(n230) );
  MAOI222D1 U178 ( .A(prm[19]), .B(n226), .C(n225), .ZN(n227) );
  NR2D1 U179 ( .A1(n243), .A2(prm[36]), .ZN(n225) );
  OAI22D1 U180 ( .A1(prm[22]), .A2(n224), .B1(prm[21]), .B2(n223), .ZN(n232)
         );
  OAI31D1 U181 ( .A1(n222), .A2(n221), .A3(n220), .B(n219), .ZN(enm[6]) );
  OAI21D1 U182 ( .A1(n218), .A2(n217), .B(n216), .ZN(n219) );
  MAOI222D1 U183 ( .A(prm[41]), .B(n96), .C(n242), .ZN(enm[11]) );
  MAOI222D1 U184 ( .A(n95), .B(prm[34]), .C(n224), .ZN(n96) );
  NR2D1 U185 ( .A1(n94), .A2(n93), .ZN(n95) );
  AOI211D1 U186 ( .A1(prm[33]), .A2(n223), .B(n92), .C(prm[32]), .ZN(n93) );
  MAOI222D1 U187 ( .A(prm[33]), .B(n91), .C(n223), .ZN(n94) );
  OAI32D1 U188 ( .A1(n89), .A2(n183), .A3(prm[36]), .B1(prm[37]), .B2(n236), 
        .ZN(n92) );
  NR2D1 U189 ( .A1(prm[31]), .A2(n226), .ZN(n89) );
  OAI211D1 U190 ( .A1(n215), .A2(n220), .B(n216), .C(n214), .ZN(enm[5]) );
  OAI21D1 U191 ( .A1(n220), .A2(n213), .B(n215), .ZN(n214) );
  CKXOR2D1 U192 ( .A1(n212), .A2(n211), .Z(n217) );
  CKXOR2D1 U193 ( .A1(n210), .A2(n209), .Z(n218) );
  AOI32D1 U194 ( .A1(n204), .A2(n203), .A3(n202), .B1(n201), .B2(n200), .ZN(
        enm[3]) );
  MAOI222D1 U195 ( .A(prm[11]), .B(n253), .C(n182), .ZN(n205) );
  MAOI222D1 U196 ( .A(prm[28]), .B(n181), .C(n180), .ZN(n182) );
  MAOI222D1 U197 ( .A(prm[9]), .B(n179), .C(n248), .ZN(n180) );
  MAOI222D1 U198 ( .A(prm[26]), .B(n178), .C(n177), .ZN(n179) );
  MAOI222D1 U199 ( .A(prm[7]), .B(n245), .C(n176), .ZN(n177) );
  NR2D1 U200 ( .A1(n175), .A2(prm[24]), .ZN(n176) );
  MAOI222D1 U201 ( .A(prm[11]), .B(n242), .C(n174), .ZN(n206) );
  MAOI222D1 U202 ( .A(prm[34]), .B(n181), .C(n173), .ZN(n174) );
  MAOI222D1 U203 ( .A(prm[9]), .B(n172), .C(n238), .ZN(n173) );
  MAOI222D1 U204 ( .A(prm[32]), .B(n178), .C(n171), .ZN(n172) );
  MAOI222D1 U205 ( .A(prm[7]), .B(n236), .C(n170), .ZN(n171) );
  NR2D1 U206 ( .A1(n175), .A2(prm[30]), .ZN(n170) );
  MAOI222D1 U207 ( .A(prm[11]), .B(n166), .C(n165), .ZN(n167) );
  MAOI222D1 U208 ( .A(prm[16]), .B(n181), .C(n164), .ZN(n165) );
  MAOI222D1 U209 ( .A(prm[9]), .B(n163), .C(n162), .ZN(n164) );
  MAOI222D1 U210 ( .A(prm[14]), .B(n161), .C(n178), .ZN(n163) );
  MAOI222D1 U211 ( .A(n160), .B(prm[7]), .C(n159), .ZN(n161) );
  NR2D1 U212 ( .A1(n175), .A2(prm[12]), .ZN(n160) );
  MAOI222D1 U213 ( .A(prm[11]), .B(n234), .C(n158), .ZN(n168) );
  OAI22D1 U214 ( .A1(prm[40]), .A2(n181), .B1(n157), .B2(n156), .ZN(n158) );
  NR2D1 U215 ( .A1(n155), .A2(n154), .ZN(n156) );
  NR2D1 U216 ( .A1(prm[39]), .A2(n153), .ZN(n154) );
  MAOI222D1 U217 ( .A(n152), .B(prm[38]), .C(n178), .ZN(n155) );
  MAOI222D1 U218 ( .A(prm[7]), .B(n226), .C(n151), .ZN(n152) );
  NR2D1 U219 ( .A1(n175), .A2(prm[36]), .ZN(n151) );
  OAI22D1 U220 ( .A1(prm[10]), .A2(n224), .B1(prm[9]), .B2(n223), .ZN(n157) );
  MAOI222D1 U221 ( .A(prm[11]), .B(n150), .C(n149), .ZN(n169) );
  MAOI222D1 U222 ( .A(prm[22]), .B(n181), .C(n148), .ZN(n149) );
  MAOI222D1 U223 ( .A(prm[9]), .B(n147), .C(n228), .ZN(n148) );
  MAOI222D1 U224 ( .A(prm[20]), .B(n178), .C(n146), .ZN(n147) );
  MAOI222D1 U225 ( .A(prm[7]), .B(n145), .C(n144), .ZN(n146) );
  NR2D1 U226 ( .A1(n175), .A2(prm[18]), .ZN(n144) );
  XNR2D1 U227 ( .A1(n261), .A2(n260), .ZN(n204) );
  MAOI222D1 U228 ( .A(prm[35]), .B(n190), .C(n253), .ZN(n261) );
  MAOI222D1 U229 ( .A(prm[28]), .B(n189), .C(n188), .ZN(n190) );
  MAOI222D1 U230 ( .A(prm[33]), .B(n248), .C(n187), .ZN(n189) );
  MAOI222D1 U231 ( .A(prm[26]), .B(n186), .C(n185), .ZN(n187) );
  MAOI222D1 U232 ( .A(prm[31]), .B(n184), .C(n245), .ZN(n186) );
  OAI21D1 U233 ( .A1(n220), .A2(n221), .B(n222), .ZN(enm[2]) );
  AO21D1 U234 ( .A1(n215), .A2(n196), .B(n213), .Z(enm[1]) );
  AOI211D1 U235 ( .A1(n142), .A2(n102), .B(n120), .C(n101), .ZN(n193) );
  NR2D1 U236 ( .A1(n142), .A2(n102), .ZN(n101) );
  NR2D1 U237 ( .A1(n100), .A2(n99), .ZN(n141) );
  NR2D1 U238 ( .A1(n98), .A2(n97), .ZN(n142) );
  AO21D1 U239 ( .A1(n122), .A2(n121), .B(n120), .Z(n197) );
  NR2D1 U240 ( .A1(n122), .A2(n121), .ZN(n120) );
  XNR2D1 U241 ( .A1(n100), .A2(n99), .ZN(n121) );
  XNR2D1 U242 ( .A1(n98), .A2(n97), .ZN(n122) );
  MAOI222D1 U243 ( .A(prm[5]), .B(n242), .C(n119), .ZN(n198) );
  MAOI222D1 U244 ( .A(prm[34]), .B(n118), .C(n117), .ZN(n119) );
  OAI21D1 U245 ( .A1(prm[3]), .A2(n238), .B(n116), .ZN(n117) );
  MAOI222D1 U246 ( .A(prm[2]), .B(n113), .C(n185), .ZN(n115) );
  MAOI222D1 U247 ( .A(prm[31]), .B(n112), .C(n111), .ZN(n113) );
  INVD1 U248 ( .I(prm[35]), .ZN(n242) );
  MAOI222D1 U249 ( .A(prm[5]), .B(n234), .C(n110), .ZN(n199) );
  MAOI222D1 U250 ( .A(prm[40]), .B(n118), .C(n109), .ZN(n110) );
  OAI21D1 U251 ( .A1(prm[3]), .A2(n223), .B(n108), .ZN(n109) );
  AOI22D1 U252 ( .A1(prm[38]), .A2(n107), .B1(n106), .B2(n105), .ZN(n108) );
  AOI22D1 U253 ( .A1(prm[2]), .A2(n104), .B1(prm[3]), .B2(n223), .ZN(n105) );
  MAOI222D1 U254 ( .A(prm[1]), .B(n226), .C(n103), .ZN(n106) );
  INR2D1 U255 ( .A1(prm[0]), .B1(prm[36]), .ZN(n103) );
  AOI21D1 U256 ( .A1(prm[3]), .A2(n223), .B(prm[2]), .ZN(n107) );
  MAOI222D1 U257 ( .A(prm[35]), .B(n127), .C(n166), .ZN(n210) );
  MAOI222D1 U258 ( .A(prm[16]), .B(n126), .C(n188), .ZN(n127) );
  MAOI222D1 U259 ( .A(prm[33]), .B(n162), .C(n125), .ZN(n126) );
  MAOI222D1 U260 ( .A(prm[14]), .B(n124), .C(n185), .ZN(n125) );
  MAOI222D1 U261 ( .A(prm[31]), .B(n123), .C(n159), .ZN(n124) );
  NR2D1 U262 ( .A1(n212), .A2(n211), .ZN(n215) );
  MAOI222D1 U263 ( .A(prm[17]), .B(n253), .C(n140), .ZN(n211) );
  MAOI222D1 U264 ( .A(prm[28]), .B(n139), .C(n138), .ZN(n140) );
  MAOI222D1 U265 ( .A(prm[15]), .B(n137), .C(n248), .ZN(n138) );
  MAOI222D1 U266 ( .A(prm[26]), .B(n136), .C(n135), .ZN(n137) );
  MAOI222D1 U267 ( .A(prm[13]), .B(n245), .C(n134), .ZN(n135) );
  NR2D1 U268 ( .A1(n133), .A2(prm[24]), .ZN(n134) );
  INVD1 U269 ( .I(prm[29]), .ZN(n253) );
  MAOI222D1 U270 ( .A(prm[17]), .B(n150), .C(n132), .ZN(n212) );
  MAOI222D1 U271 ( .A(prm[22]), .B(n139), .C(n131), .ZN(n132) );
  MAOI222D1 U272 ( .A(n130), .B(prm[15]), .C(n228), .ZN(n131) );
  MAOI222D1 U273 ( .A(prm[20]), .B(n129), .C(n136), .ZN(n130) );
  MAOI222D1 U274 ( .A(prm[13]), .B(n145), .C(n128), .ZN(n129) );
  NR2D1 U275 ( .A1(n133), .A2(prm[18]), .ZN(n128) );
  FA1D0 U276 ( .A(n169), .B(n168), .CI(n167), .CO(n201), .S(n207) );
  MUX2ND0 U277 ( .I0(n195), .I1(n194), .S(n193), .ZN(n213) );
  FA1D0 U278 ( .A(n199), .B(n198), .CI(n197), .CO(n194), .S(n222) );
  FA1D0 U279 ( .A(n207), .B(n206), .CI(n205), .CO(n200), .S(n208) );
  FA1D0 U280 ( .A(n257), .B(n256), .CI(n255), .CO(n254), .S(n258) );
endmodule

