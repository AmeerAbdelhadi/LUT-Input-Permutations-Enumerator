
module enumerate ( prm, enm );
  input [35:0] prm;
  output [8:0] enm;
  wire   n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165;

  CKND2D0 U38 ( .A1(n165), .A2(n164), .ZN(enm[7]) );
  CKND2D0 U39 ( .A1(n161), .A2(n160), .ZN(n165) );
  CKND0 U40 ( .I(n80), .ZN(n160) );
  CKND0 U41 ( .I(n81), .ZN(n161) );
  CKND0 U42 ( .I(n159), .ZN(enm[5]) );
  CKND0 U43 ( .I(n155), .ZN(enm[4]) );
  CKND0 U44 ( .I(prm[12]), .ZN(n144) );
  CKND0 U45 ( .I(prm[14]), .ZN(n148) );
  CKND0 U46 ( .I(prm[34]), .ZN(n35) );
  CKND0 U47 ( .I(prm[32]), .ZN(n32) );
  CKND0 U48 ( .I(prm[24]), .ZN(n30) );
  CKND2D0 U49 ( .A1(n124), .A2(n123), .ZN(n122) );
  CKND2D0 U50 ( .A1(n127), .A2(n126), .ZN(n125) );
  CKND2D0 U51 ( .A1(n120), .A2(n121), .ZN(n123) );
  CKND0 U52 ( .I(n114), .ZN(n115) );
  CKND0 U53 ( .I(prm[16]), .ZN(n152) );
  CKND0 U54 ( .I(prm[22]), .ZN(n104) );
  CKND0 U55 ( .I(prm[20]), .ZN(n100) );
  CKND2D0 U56 ( .A1(prm[6]), .A2(n97), .ZN(n99) );
  CKND0 U57 ( .I(prm[18]), .ZN(n97) );
  CKND0 U58 ( .I(prm[6]), .ZN(n107) );
  CKND0 U59 ( .I(prm[8]), .ZN(n111) );
  CKND0 U60 ( .I(prm[10]), .ZN(n95) );
  CKND0 U61 ( .I(n85), .ZN(enm[1]) );
  CKND0 U62 ( .I(prm[21]), .ZN(n149) );
  CKND0 U63 ( .I(prm[19]), .ZN(n146) );
  CKND0 U64 ( .I(prm[23]), .ZN(n154) );
  CKND0 U65 ( .I(prm[27]), .ZN(n139) );
  CKND0 U66 ( .I(prm[25]), .ZN(n137) );
  CKND0 U67 ( .I(prm[9]), .ZN(n103) );
  CKND0 U68 ( .I(prm[7]), .ZN(n98) );
  CKND0 U69 ( .I(prm[11]), .ZN(n117) );
  CKND0 U70 ( .I(prm[33]), .ZN(n131) );
  CKND0 U71 ( .I(prm[31]), .ZN(n129) );
  CKND0 U72 ( .I(prm[35]), .ZN(n135) );
  CKND0 U73 ( .I(prm[15]), .ZN(n112) );
  CKND0 U74 ( .I(prm[0]), .ZN(n69) );
  CKND0 U75 ( .I(prm[13]), .ZN(n108) );
  CKND0 U76 ( .I(prm[2]), .ZN(n72) );
  CKND0 U77 ( .I(prm[4]), .ZN(n75) );
  CKND0 U78 ( .I(prm[17]), .ZN(n53) );
  AOI32D1 U79 ( .A1(n164), .A2(n160), .A3(n161), .B1(n81), .B2(n80), .ZN(
        enm[0]) );
  XNR2D1 U80 ( .A1(n163), .A2(n162), .ZN(n164) );
  OAI21D1 U81 ( .A1(n163), .A2(n162), .B(n165), .ZN(enm[6]) );
  MAOI222D1 U82 ( .A(prm[23]), .B(n143), .C(n47), .ZN(n162) );
  MAOI222D1 U83 ( .A(prm[28]), .B(n104), .C(n46), .ZN(n47) );
  MAOI222D1 U84 ( .A(n45), .B(prm[21]), .C(n139), .ZN(n46) );
  MAOI222D1 U85 ( .A(prm[26]), .B(n44), .C(n100), .ZN(n45) );
  MAOI222D1 U86 ( .A(prm[19]), .B(n137), .C(n43), .ZN(n44) );
  NR2D1 U87 ( .A1(n97), .A2(prm[24]), .ZN(n43) );
  MAOI222D1 U88 ( .A(prm[23]), .B(n135), .C(n42), .ZN(n163) );
  MAOI222D1 U89 ( .A(prm[34]), .B(n104), .C(n41), .ZN(n42) );
  MAOI222D1 U90 ( .A(prm[21]), .B(n40), .C(n131), .ZN(n41) );
  MAOI222D1 U91 ( .A(prm[32]), .B(n100), .C(n39), .ZN(n40) );
  MAOI222D1 U92 ( .A(prm[19]), .B(n129), .C(n38), .ZN(n39) );
  NR2D1 U93 ( .A1(n97), .A2(prm[30]), .ZN(n38) );
  MAOI222D1 U94 ( .A(prm[17]), .B(n154), .C(n153), .ZN(n156) );
  MAOI222D1 U95 ( .A(prm[22]), .B(n152), .C(n151), .ZN(n153) );
  MAOI222D1 U96 ( .A(prm[15]), .B(n150), .C(n149), .ZN(n151) );
  MAOI222D1 U97 ( .A(prm[20]), .B(n148), .C(n147), .ZN(n150) );
  MAOI222D1 U98 ( .A(prm[13]), .B(n146), .C(n145), .ZN(n147) );
  NR2D1 U99 ( .A1(n144), .A2(prm[18]), .ZN(n145) );
  MAOI222D1 U100 ( .A(prm[17]), .B(n143), .C(n142), .ZN(n157) );
  MAOI222D1 U101 ( .A(prm[28]), .B(n152), .C(n141), .ZN(n142) );
  MAOI222D1 U102 ( .A(prm[15]), .B(n140), .C(n139), .ZN(n141) );
  MAOI222D1 U103 ( .A(prm[26]), .B(n148), .C(n138), .ZN(n140) );
  MAOI222D1 U104 ( .A(prm[13]), .B(n137), .C(n136), .ZN(n138) );
  NR2D1 U105 ( .A1(n144), .A2(prm[24]), .ZN(n136) );
  MAOI222D1 U106 ( .A(prm[17]), .B(n135), .C(n134), .ZN(n158) );
  MAOI222D1 U107 ( .A(prm[34]), .B(n152), .C(n133), .ZN(n134) );
  MAOI222D1 U108 ( .A(prm[15]), .B(n132), .C(n131), .ZN(n133) );
  MAOI222D1 U109 ( .A(prm[32]), .B(n148), .C(n130), .ZN(n132) );
  MAOI222D1 U110 ( .A(prm[13]), .B(n129), .C(n128), .ZN(n130) );
  NR2D1 U111 ( .A1(n144), .A2(prm[30]), .ZN(n128) );
  MAOI222D1 U112 ( .A(prm[35]), .B(n37), .C(n143), .ZN(enm[8]) );
  MAOI222D1 U113 ( .A(prm[28]), .B(n36), .C(n35), .ZN(n37) );
  MAOI222D1 U114 ( .A(prm[33]), .B(n139), .C(n34), .ZN(n36) );
  MAOI222D1 U115 ( .A(prm[26]), .B(n33), .C(n32), .ZN(n34) );
  OAI32D1 U116 ( .A1(n31), .A2(n30), .A3(prm[30]), .B1(prm[31]), .B2(n137), 
        .ZN(n33) );
  NR2D1 U117 ( .A1(prm[25]), .A2(n129), .ZN(n31) );
  OA21D1 U118 ( .A1(n127), .A2(n126), .B(n125), .Z(enm[3]) );
  OAI211D1 U119 ( .A1(n124), .A2(n123), .B(n125), .C(n122), .ZN(enm[2]) );
  CKXOR2D1 U120 ( .A1(n121), .A2(n120), .Z(n126) );
  CKXOR2D1 U121 ( .A1(n119), .A2(n118), .Z(n127) );
  MAOI222D1 U122 ( .A(n117), .B(prm[17]), .C(n116), .ZN(n121) );
  MAOI222D1 U123 ( .A(n152), .B(prm[10]), .C(n115), .ZN(n116) );
  MAOI222D1 U124 ( .A(prm[9]), .B(n113), .C(n112), .ZN(n114) );
  MAOI222D1 U125 ( .A(prm[14]), .B(n111), .C(n110), .ZN(n113) );
  MAOI222D1 U126 ( .A(prm[7]), .B(n109), .C(n108), .ZN(n110) );
  NR2D1 U127 ( .A1(prm[12]), .A2(n107), .ZN(n109) );
  MAOI222D1 U128 ( .A(prm[23]), .B(n106), .C(n117), .ZN(n120) );
  MAOI222D1 U129 ( .A(prm[10]), .B(n105), .C(n104), .ZN(n106) );
  MAOI222D1 U130 ( .A(prm[21]), .B(n103), .C(n102), .ZN(n105) );
  MAOI222D1 U131 ( .A(prm[8]), .B(n101), .C(n100), .ZN(n102) );
  MAOI222D1 U132 ( .A(prm[19]), .B(n99), .C(n98), .ZN(n101) );
  NR2D1 U133 ( .A1(n119), .A2(n118), .ZN(n124) );
  MAOI222D1 U134 ( .A(prm[11]), .B(n135), .C(n96), .ZN(n118) );
  MAOI222D1 U135 ( .A(prm[34]), .B(n95), .C(n94), .ZN(n96) );
  MAOI222D1 U136 ( .A(prm[9]), .B(n93), .C(n131), .ZN(n94) );
  MAOI222D1 U137 ( .A(prm[32]), .B(n111), .C(n92), .ZN(n93) );
  MAOI222D1 U138 ( .A(prm[7]), .B(n129), .C(n91), .ZN(n92) );
  NR2D1 U139 ( .A1(n107), .A2(prm[30]), .ZN(n91) );
  MAOI222D1 U140 ( .A(prm[11]), .B(n143), .C(n90), .ZN(n119) );
  MAOI222D1 U141 ( .A(prm[28]), .B(n95), .C(n89), .ZN(n90) );
  MAOI222D1 U142 ( .A(prm[9]), .B(n88), .C(n139), .ZN(n89) );
  MAOI222D1 U143 ( .A(prm[26]), .B(n111), .C(n87), .ZN(n88) );
  MAOI222D1 U144 ( .A(prm[7]), .B(n137), .C(n86), .ZN(n87) );
  NR2D1 U145 ( .A1(n107), .A2(prm[24]), .ZN(n86) );
  MAOI222D1 U146 ( .A(prm[5]), .B(n154), .C(n76), .ZN(n82) );
  MAOI222D1 U147 ( .A(prm[22]), .B(n75), .C(n74), .ZN(n76) );
  MAOI222D1 U148 ( .A(prm[3]), .B(n73), .C(n149), .ZN(n74) );
  MAOI222D1 U149 ( .A(prm[20]), .B(n72), .C(n71), .ZN(n73) );
  MAOI222D1 U150 ( .A(prm[1]), .B(n146), .C(n70), .ZN(n71) );
  NR2D1 U151 ( .A1(n69), .A2(prm[18]), .ZN(n70) );
  MAOI222D1 U152 ( .A(prm[5]), .B(n143), .C(n68), .ZN(n83) );
  MAOI222D1 U153 ( .A(prm[28]), .B(n75), .C(n67), .ZN(n68) );
  MAOI222D1 U154 ( .A(prm[3]), .B(n66), .C(n139), .ZN(n67) );
  MAOI222D1 U155 ( .A(prm[26]), .B(n72), .C(n65), .ZN(n66) );
  MAOI222D1 U156 ( .A(prm[1]), .B(n137), .C(n64), .ZN(n65) );
  NR2D1 U157 ( .A1(n69), .A2(prm[24]), .ZN(n64) );
  INVD1 U158 ( .I(prm[29]), .ZN(n143) );
  MAOI222D1 U159 ( .A(prm[5]), .B(n117), .C(n63), .ZN(n77) );
  MAOI222D1 U160 ( .A(prm[10]), .B(n75), .C(n62), .ZN(n63) );
  MAOI222D1 U161 ( .A(prm[3]), .B(n61), .C(n103), .ZN(n62) );
  MAOI222D1 U162 ( .A(prm[8]), .B(n72), .C(n60), .ZN(n61) );
  MAOI222D1 U163 ( .A(prm[1]), .B(n98), .C(n59), .ZN(n60) );
  NR2D1 U164 ( .A1(n69), .A2(prm[6]), .ZN(n59) );
  MAOI222D1 U165 ( .A(prm[5]), .B(n135), .C(n58), .ZN(n78) );
  MAOI222D1 U166 ( .A(prm[34]), .B(n75), .C(n57), .ZN(n58) );
  MAOI222D1 U167 ( .A(prm[3]), .B(n56), .C(n131), .ZN(n57) );
  MAOI222D1 U168 ( .A(prm[32]), .B(n72), .C(n55), .ZN(n56) );
  MAOI222D1 U169 ( .A(prm[1]), .B(n129), .C(n54), .ZN(n55) );
  NR2D1 U170 ( .A1(n69), .A2(prm[30]), .ZN(n54) );
  MAOI222D1 U171 ( .A(prm[5]), .B(n53), .C(n52), .ZN(n79) );
  MAOI222D1 U172 ( .A(prm[16]), .B(n75), .C(n51), .ZN(n52) );
  MAOI222D1 U173 ( .A(prm[3]), .B(n50), .C(n112), .ZN(n51) );
  MAOI222D1 U174 ( .A(prm[14]), .B(n72), .C(n49), .ZN(n50) );
  MAOI222D1 U175 ( .A(prm[1]), .B(n108), .C(n48), .ZN(n49) );
  NR2D1 U176 ( .A1(n69), .A2(prm[12]), .ZN(n48) );
  FA1D0 U177 ( .A(n79), .B(n78), .CI(n77), .CO(n81), .S(n84) );
  FA1D0 U178 ( .A(n84), .B(n83), .CI(n82), .CO(n80), .S(n85) );
  FA1D0 U179 ( .A(n158), .B(n157), .CI(n156), .CO(n155), .S(n159) );
endmodule

